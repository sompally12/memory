module tb;
endmodule
