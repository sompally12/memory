interface mem_if;
endinterface
